module fa(
input a,b,c,output s,y);
assign {y,s}=a+b+c;
endmodule